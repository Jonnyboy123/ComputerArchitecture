module PCArith(PC, Add, InstructionCache);

	input PC, Add;
	output InstructionCache;
	
	 
endmodule 