module DataCache(Address, WriteData, ReadData, DataMem);

	input Address, WriteData;
	output ReadData, DataMem;
	
endmodule 