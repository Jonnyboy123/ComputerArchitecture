module OperandPrep(ReadReg1, ReadReg2, WriteReg, WriteData, ReadData1, ReadData2);

	input ReadReg1, ReadReg2, WriteReg, WriteData;
	output ReadData1, ReadData2;
	
endmodule 