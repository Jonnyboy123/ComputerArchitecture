module instruction_cache(read_address, instruction, instructionmem);

		input read_address;
		output instruction, instructionmem;
		
endmodule 